-------------------------------------------------------
--! @file
--! @author Julian Mendez <julian.mendez@cern.ch> (CERN - EP-ESE-BE)
--! @version 6.0
--! @brief GBT-FPGA IP - Rx Gearbox
-------------------------------------------------------

--! Include the IEEE VHDL standard library
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Include the GBT-FPGA specific packages
use work.gbt_bank_package.all;
use work.vendor_specific_gbt_bank_package.all;

--! @brief GBT_rx_gearbox - Rx Gearbox
--! @details 
--! The Rx gearbox module is used to ensure the MGT to Datapath clock domain
--! crossing. It takes the 20/40bit words in input and generates an 120bit
--! word every 3/6 clock cycle.
entity gbt_rx_gearbox is
  generic ( 
    RX_OPTIMIZATION           : integer range 0 to 1 := STANDARD               --! RX_OPTIMIZATION: Latency mode for the Rx path (STANDARD or LATENCY_OPTIMIZED)
  );
  port (  
    --================--
    -- Reset & Clocks --
    --================--    
    RX_RESET_I                : in  std_logic;                                  --! Reset the Rx gearbox (Asynchronous)
    RX_WORDCLK_I              : in  std_logic;                                  --! Recovered clock from data generated by the transceiver
    RX_FRAMECLK_I             : in  std_logic;
	 RX_CLKEN_i                : in  std_logic;
	 RX_CLKEN_o                : out  std_logic;
    --==============--
    -- Control      --
    --==============--
    RX_HEADERFLAG_i           : in  std_logic;                                  --! Pulsed during the clock cycle of the header
    READY_O                   : out std_logic;
	 
    --==============--
    -- Word & Frame --
    --==============--      
    RX_WORD_I                 : in  std_logic_vector(WORD_WIDTH-1 downto 0);    --! 20/40bit word from the transceiver
    RX_FRAME_O                : out std_logic_vector(119 downto 0)              --! 120bit aligned to be decoded
      
   );   
end gbt_rx_gearbox;

--! @brief GBT_rx_gearbox architecture - Rx Gearbox
--! @details Two gearboxes can be implemented to ensure the clock domain crossing:
--!     * *Standard mode*: The standard mode is based on a device specific IP in order to simplify the clock domain crossing. Nevertheless, this method increases the latency and might be not fix depending on the manufacturer.
--!     * *Latency Optimized*: The latency optimized mode is based on a single register where the word is saved before being pushed in output at the header flag clock cycle. 
architecture structural of gbt_rx_gearbox is
begin
   
   --==================================== User Logic =====================================--
   
    --! Instiation of the Rx gearbox (Standard mode)
    rxGearboxStd_gen: if RX_OPTIMIZATION = STANDARD generate
      rxGearboxStd: entity work.gbt_rx_gearbox_std
         port map (           
             RX_RESET_I                                => RX_RESET_I,
      
             RX_WORDCLK_I                              => RX_WORDCLK_I,
             RX_FRAMECLK_I                             => RX_FRAMECLK_I,
				 RX_CLKEN_i                                => RX_CLKEN_i,
             RX_CLKEN_o                                => RX_CLKEN_o,
				 
             READY_O                                   => READY_O,
             Rx_HEADERFLAG_i                           => Rx_HEADERFLAG_i,
      
             RX_WORD_I                                 => RX_WORD_I,
             RX_FRAME_O                                => RX_FRAME_O    
         );     
    end generate;   
   
    --! Instiation of the Rx gearbox (Latency optimized mode)
    rxGearboxLatOpt_gen: if RX_OPTIMIZATION = LATENCY_OPTIMIZED generate   
      rxGearboxLatOpt: entity work.gbt_rx_gearbox_latopt
        port map (   
          RX_RESET_I                  => RX_RESET_I,
          RX_WORDCLK_I                => RX_WORDCLK_I,
			 RX_FRAMECLK_I               => RX_FRAMECLK_I,
			 RX_CLKEN_i                  => RX_CLKEN_i,
          RX_HEADERFLAG_i             => RX_HEADERFLAG_i,
			 RX_CLKEN_o                  => RX_CLKEN_o,
			 READY_O                     => READY_O,
          RX_WORD_I                   => RX_WORD_I,
          RX_FRAME_O                  => RX_FRAME_O
        );
   end generate;
   
   --=====================================================================================--   
end structural;
--=================================================================================================--
--#################################################################################################--
--=================================================================================================--